* rc_common
.param
+ tc1rsn=1.422e-3
+ tc2rsn=6.569e-7
+ tc1rsp=1.259e-3
+ tc2rsp=2.204e-6
+ tc1rsn_h=1.405e-3
+ tc2rsn_h=4.233e-7
+ tc1rsp_h=1.369e-3
+ tc2rsp_h=1.476e-6
+ tc1rsnw=1.483e-3
+ tc2rsnw=7.824e-6
+ tc1rsgpu=8.916e-4
+ tc2rsgpu=8.443e-7
+ nfom_dw=0.017u
+ pfom_dw=0.004u
+ poly_dw=-0.056u
+ li_dw=0.017u
+ m1_dw=-0.039u
+ m2_dw=-0.039u
+ m3_dw=-0.025u
+ m4_dw=-0.025u
+ m5_dw=-0.09u
+ rdl_dw=0.0u
