* C4M.Sky130 global per device corner lib file

.lib logic_tt
.include "C4M.Sky130_logic_tt_model.spice"
.endl logic_tt
.lib logic_ff
.include "C4M.Sky130_logic_ff_model.spice"
.endl logic_ff
.lib logic_ss
.include "C4M.Sky130_logic_ss_model.spice"
.endl logic_ss
.lib logic_fs
.include "C4M.Sky130_logic_fs_model.spice"
.endl logic_fs
.lib logic_sf
.include "C4M.Sky130_logic_sf_model.spice"
.endl logic_sf
.lib io_tt
.include "C4M.Sky130_io_tt_model.spice"
.endl io_tt
.lib io_ff
.include "C4M.Sky130_io_ff_model.spice"
.endl io_ff
.lib io_ss
.include "C4M.Sky130_io_ss_model.spice"
.endl io_ss
.lib io_fs
.include "C4M.Sky130_io_fs_model.spice"
.endl io_fs
.lib io_sf
.include "C4M.Sky130_io_sf_model.spice"
.endl io_sf
.lib diode_tt
.include "C4M.Sky130_diode_tt_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl diode_tt
.lib diode_ff
.include "C4M.Sky130_diode_ff_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl diode_ff
.lib diode_ss
.include "C4M.Sky130_diode_ss_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl diode_ss
.lib diode_fs
.include "C4M.Sky130_diode_fs_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl diode_fs
.lib diode_sf
.include "C4M.Sky130_diode_sf_params.spice"
.include "C4M.Sky130_diode_model.spice"
.endl diode_sf
.lib pnp_t
.include "C4M.Sky130_pnp_t_params.spice"
.include "C4M.Sky130_pnp_model.spice"
.endl npn_t
.lib pnp_f
.include "C4M.Sky130_pnp_f_params.spice"
.include "C4M.Sky130_pnp_model.spice"
.endl npn_f
.lib pnp_s
.include "C4M.Sky130_pnp_s_params.spice"
.include "C4M.Sky130_pnp_model.spice"
.endl npn_s
.lib npn_t
.include "C4M.Sky130_npn_t_params.spice"
.include "C4M.Sky130_npn_model.spice"
.endl npn_t
.lib npn_f
.include "C4M.Sky130_npn_f_params.spice"
.include "C4M.Sky130_npn_model.spice"
.endl npn_f
.lib npn_s
.include "C4M.Sky130_npn_s_params.spice"
.include "C4M.Sky130_npn_model.spice"
.endl npn_s
.lib rc_tt
.include "C4M.Sky130_rc_tt_params.spice"
.include "C4M.Sky130_rc_common_params.spice"
.include "C4M.Sky130_rc_model.spice"
.endl rc_tt
.lib rc_ll
.include "C4M.Sky130_rc_ll_params.spice"
.include "C4M.Sky130_rc_common_params.spice"
.include "C4M.Sky130_rc_model.spice"
.endl rc_ll
.lib rc_hh
.include "C4M.Sky130_rc_hh_params.spice"
.include "C4M.Sky130_rc_common_params.spice"
.include "C4M.Sky130_rc_model.spice"
.endl rc_hh
.lib rc_lh
.include "C4M.Sky130_rc_lh_params.spice"
.include "C4M.Sky130_rc_common_params.spice"
.include "C4M.Sky130_rc_model.spice"
.endl rc_lh
.lib rc_hl
.include "C4M.Sky130_rc_hl_params.spice"
.include "C4M.Sky130_rc_common_params.spice"
.include "C4M.Sky130_rc_model.spice"
.endl rc_hl
