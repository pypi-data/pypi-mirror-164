* rc_tt
.param
+ tol_nfom=0
+ tol_pfom=0
+ tol_nw=0.0
+ tol_poly=0.0
+ tol_li=0.0
+ tol_m1=0.0
+ tol_m2=0.0
+ tol_m3=0.0
+ tol_m4=0.0
+ tol_m5=0.0
+ tol_rdl=0.0
+ rdn=120
+ rdp=197
+ rdn_hv=114
+ rdp_hv=191
+ rp1=48.2
+ rnw=1700
+ rl1=12.2
+ rm1=0.125
+ rm2=0.125
+ rm3=0.047
+ rm4=0.047
+ rm5=0.0285
+ rrdl=0.005
